* nupa

* (exec-spice "ngspice %s")
* (compile "cd ../w32 && LC_ALL=eC make -k")
*
* check ?: assoziativity

.param foo_1001 = '3>2 ? 42 : 3>2 ? 41 : 40'
.param foo_1002 = '3>2 ? 42 : 3<2 ? 41 : 40'
.param foo_1003 = '3<2 ? 42 : 3>2 ? 41 : 40'
.param foo_1004 = '3<2 ? 42 : 3<2 ? 41 : 40'

v1001  1001 0  'foo_1001'
v1002  1002 0  'foo_1002'
v1003  1003 0  'foo_1003'
v1004  1004 0  'foo_1004'

.control

define mismatch(a,b,err) abs(a-b)>err

op

let baz_1001 = (3 gt 2 ? 42 : 3 gt 2 ? 41 : 40)
let baz_1002 = (3 gt 2 ? 42 : 3 lt 2 ? 41 : 40)
let baz_1003 = (3 lt 2 ? 42 : 3 gt 2 ? 41 : 40)
let baz_1004 = (3 lt 2 ? 42 : 3 lt 2 ? 41 : 40)

print all

if mismatch(v(1001), 42, 1e-9)
  echo "ERROR, mismatch 1001"
end

if mismatch(v(1002), 42, 1e-9)
  echo "ERROR, mismatch 1002"
end

if mismatch(v(1003), 41, 1e-9)
  echo "ERROR, mismatch 1003"
end

if mismatch(v(1004), 40, 1e-9)
  echo "ERROR, mismatch 1004"
end

quit 1

.endc
