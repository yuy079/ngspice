check current transfer function
* (compile "../w32/src/ngspice tf-3.cir" t)

iin  0 1  DC=8mA
r1   1 2  100
d1   2 0  Dmod

.model Dmod D(IS=10f)

.control

let vt = boltz * (27.0 - kelvin) / echarge

op 

let rd = const.vt / @d1[id]

let gold_Zout = rd
let gold_Zin  = @r1[resistance] + rd
let gold_tf   = rd

tf v(2) iin
print all

define relerr(y,gold) (y/gold - 1)

echo "--"

print relerr(transfer_function, op1.gold_tf)
print relerr(iin#input_impedance, op1.gold_Zin)
print relerr(output_impedance_at_v(2), op1.gold_Zout)

.endc

.end
